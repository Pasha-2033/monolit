`ifndef STD_UTILS
	`include "utils.sv"
`endif
`define STD_IO
`include "io/SPI.sv"