module ALU #(
	parameter word_width
) (
	input wire	[word_width - 1:0]	A,
	input wire	[word_width - 1:0]	B,
	output wire	[word_width - 1:0]	R
);

endmodule