`include "utils.sv"
`include "tree_decoder.sv"
`include "CLAA.sv"
`include "CSA_S.sv"
`include "fast_comparator.sv"
`include "polyshift_r.sv"
`include "polyshift_l.sv"
`include "RCA_M.sv"
`include "screening_by_junior.sv"
`include "screening_by_senior.sv"
`timescale 1ps/1ps
module utils_tb;
task_tree_decoder #(.OUTPUT_WIDTH(12)) td();
task_CLAA #(.WORD_WIDTH(16)) claa();
task_CSA_S #(.WORD_WIDTH(12), .UNIT_WIDTH(5)) csa_s();
task_fast_comparator #(.WORD_WIDTH(7)) fc();
task_polyshift_r #(.WORD_WIDTH(8)) psr();
task_polyshift_l #(.WORD_WIDTH(8)) psl();
task_RCA_M #(.WORD_WIDTH(16)) rca_m();
task_screening_by_junior #(.WORD_WIDTH(8)) sbj();
task_screening_by_senior #(.WORD_WIDTH(8)) sbs();
initial begin
	$display("_tree_decoder task:");
	td.run(0);
	td.run(1);
	td.run(2);
	td.run(10);
	td.run(11);
	$display("CLAA task:");
	repeat (10) begin
		claa.run($urandom, $urandom);
	end
	$display("CSA_S task:");
	repeat (10) begin
		csa_s.run($urandom, $urandom);
	end
	$display("fast_comparator task:");
	fc.run(2, 1);
	fc.run(1, 2);
	fc.run(15, 14);
	fc.run(12, 13);
	fc.run(11, 11);
	fc.run(20, 78);
	fc.run(123, 100);
	$display("polyshift_r task:");
	psr.run(8'b11001100, 7'b0101010);
	$display("polyshift_l task:");
	psl.run(8'b00110011, 7'b1010101);
	$display("RCA_M task:");
	repeat (10) begin
		rca_m.run($urandom, $urandom);
	end
	$display("screening_by_junior task:");
	repeat (10) begin
		sbj.run($urandom);
	end
	$display("screening_by_senior task:");
	repeat (10) begin
		sbs.run($urandom);
	end
end
endmodule